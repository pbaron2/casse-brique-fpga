-- Niosballe.vhd

-- Generated using ACDS version 18.0 614

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Niosballe is
	port (
		adr_brique_export   : out   std_logic_vector(8 downto 0);                     --   adr_brique.export
		brique_morte_export : in    std_logic                     := '0';             -- brique_morte.export
		clk_clk             : in    std_logic                     := '0';             --          clk.clk
		en_export           : in    std_logic                     := '0';             --           en.export
		en_nios_export      : out   std_logic;                                        --      en_nios.export
		fincalcul_export    : out   std_logic;                                        --    fincalcul.export
		perdu_export        : out   std_logic;                                        --        perdu.export
		pos_raquette_export : in    std_logic_vector(10 downto 0) := (others => '0'); -- pos_raquette.export
		reset_reset_n       : in    std_logic                     := '0';             --        reset.reset_n
		sram_de2_ADDR       : out   std_logic_vector(17 downto 0);                    --     sram_de2.ADDR
		sram_de2_DQ         : inout std_logic_vector(15 downto 0) := (others => '0'); --             .DQ
		sram_de2_WE_N       : out   std_logic;                                        --             .WE_N
		sram_de2_OE_N       : out   std_logic;                                        --             .OE_N
		sram_de2_UB_N       : out   std_logic;                                        --             .UB_N
		sram_de2_LB_N       : out   std_logic;                                        --             .LB_N
		sram_de2_CE_N       : out   std_logic;                                        --             .CE_N
		x_position_export   : out   std_logic_vector(10 downto 0);                    --   x_position.export
		y_position_export   : out   std_logic_vector(10 downto 0)                     --   y_position.export
	);
end entity Niosballe;

architecture rtl of Niosballe is
	component SRAM_DE2 is
		port (
			clk               : in    std_logic                     := 'X';             -- clk
			reset_n           : in    std_logic                     := 'X';             -- reset_n
			avs_s0_readdata   : out   std_logic_vector(15 downto 0);                    -- readdata
			avs_s0_writedata  : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			avs_s0_address    : in    std_logic_vector(17 downto 0) := (others => 'X'); -- address
			avs_s0_write      : in    std_logic                     := 'X';             -- write
			avs_s0_read       : in    std_logic                     := 'X';             -- read
			avs_s0_byteenable : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			coe_SRAM_ADDR     : out   std_logic_vector(17 downto 0);                    -- export
			coe_SRAM_DQ       : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			coe_SRAM_WE_N     : out   std_logic;                                        -- export
			coe_SRAM_OE_N     : out   std_logic;                                        -- export
			coe_SRAM_UB_N     : out   std_logic;                                        -- export
			coe_SRAM_LB_N     : out   std_logic;                                        -- export
			coe_SRAM_CE_N     : out   std_logic                                         -- export
		);
	end component SRAM_DE2;

	component Niosballe_adr_brique is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(8 downto 0)                      -- export
		);
	end component Niosballe_adr_brique;

	component Niosballe_brique_morte is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic                     := 'X'              -- export
		);
	end component Niosballe_brique_morte;

	component Niosballe_en_nios is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic                                         -- export
		);
	end component Niosballe_en_nios;

	component Niosballe_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component Niosballe_jtag_uart_0;

	component Niosballe_nios2_gen2_0 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(20 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(20 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component Niosballe_nios2_gen2_0;

	component Niosballe_pos_raquette is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(10 downto 0) := (others => 'X')  -- export
		);
	end component Niosballe_pos_raquette;

	component Niosballe_x_position is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(10 downto 0)                     -- export
		);
	end component Niosballe_x_position;

	component Niosballe_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                  : in  std_logic                     := 'X';             -- clk
			nios2_gen2_0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			nios2_gen2_0_data_master_address               : in  std_logic_vector(20 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_data_master_waitrequest           : out std_logic;                                        -- waitrequest
			nios2_gen2_0_data_master_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_gen2_0_data_master_read                  : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_data_master_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_gen2_0_data_master_readdatavalid         : out std_logic;                                        -- readdatavalid
			nios2_gen2_0_data_master_write                 : in  std_logic                     := 'X';             -- write
			nios2_gen2_0_data_master_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_gen2_0_data_master_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			nios2_gen2_0_instruction_master_address        : in  std_logic_vector(20 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_instruction_master_waitrequest    : out std_logic;                                        -- waitrequest
			nios2_gen2_0_instruction_master_read           : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_instruction_master_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_gen2_0_instruction_master_readdatavalid  : out std_logic;                                        -- readdatavalid
			adr_brique_s1_address                          : out std_logic_vector(1 downto 0);                     -- address
			adr_brique_s1_write                            : out std_logic;                                        -- write
			adr_brique_s1_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			adr_brique_s1_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			adr_brique_s1_chipselect                       : out std_logic;                                        -- chipselect
			brique_morte_s1_address                        : out std_logic_vector(1 downto 0);                     -- address
			brique_morte_s1_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			en_s1_address                                  : out std_logic_vector(1 downto 0);                     -- address
			en_s1_readdata                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			en_nios_s1_address                             : out std_logic_vector(1 downto 0);                     -- address
			en_nios_s1_write                               : out std_logic;                                        -- write
			en_nios_s1_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			en_nios_s1_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			en_nios_s1_chipselect                          : out std_logic;                                        -- chipselect
			fincalcul_s1_address                           : out std_logic_vector(1 downto 0);                     -- address
			fincalcul_s1_write                             : out std_logic;                                        -- write
			fincalcul_s1_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			fincalcul_s1_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			fincalcul_s1_chipselect                        : out std_logic;                                        -- chipselect
			jtag_uart_0_avalon_jtag_slave_address          : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_0_avalon_jtag_slave_write            : out std_logic;                                        -- write
			jtag_uart_0_avalon_jtag_slave_read             : out std_logic;                                        -- read
			jtag_uart_0_avalon_jtag_slave_readdata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_writedata        : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest      : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect       : out std_logic;                                        -- chipselect
			nios2_gen2_0_debug_mem_slave_address           : out std_logic_vector(8 downto 0);                     -- address
			nios2_gen2_0_debug_mem_slave_write             : out std_logic;                                        -- write
			nios2_gen2_0_debug_mem_slave_read              : out std_logic;                                        -- read
			nios2_gen2_0_debug_mem_slave_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_gen2_0_debug_mem_slave_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_gen2_0_debug_mem_slave_byteenable        : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess       : out std_logic;                                        -- debugaccess
			perdu_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			perdu_s1_write                                 : out std_logic;                                        -- write
			perdu_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			perdu_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			perdu_s1_chipselect                            : out std_logic;                                        -- chipselect
			pos_raquette_s1_address                        : out std_logic_vector(1 downto 0);                     -- address
			pos_raquette_s1_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			SRAM_DE2_0_s0_address                          : out std_logic_vector(17 downto 0);                    -- address
			SRAM_DE2_0_s0_write                            : out std_logic;                                        -- write
			SRAM_DE2_0_s0_read                             : out std_logic;                                        -- read
			SRAM_DE2_0_s0_readdata                         : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			SRAM_DE2_0_s0_writedata                        : out std_logic_vector(15 downto 0);                    -- writedata
			SRAM_DE2_0_s0_byteenable                       : out std_logic_vector(1 downto 0);                     -- byteenable
			x_position_s1_address                          : out std_logic_vector(1 downto 0);                     -- address
			x_position_s1_write                            : out std_logic;                                        -- write
			x_position_s1_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			x_position_s1_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			x_position_s1_chipselect                       : out std_logic;                                        -- chipselect
			y_position_s1_address                          : out std_logic_vector(1 downto 0);                     -- address
			y_position_s1_write                            : out std_logic;                                        -- write
			y_position_s1_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			y_position_s1_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			y_position_s1_chipselect                       : out std_logic                                         -- chipselect
		);
	end component Niosballe_mm_interconnect_0;

	component Niosballe_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component Niosballe_irq_mapper;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal nios2_gen2_0_data_master_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	signal nios2_gen2_0_data_master_waitrequest                            : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	signal nios2_gen2_0_data_master_debugaccess                            : std_logic;                     -- nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	signal nios2_gen2_0_data_master_address                                : std_logic_vector(20 downto 0); -- nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	signal nios2_gen2_0_data_master_byteenable                             : std_logic_vector(3 downto 0);  -- nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	signal nios2_gen2_0_data_master_read                                   : std_logic;                     -- nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	signal nios2_gen2_0_data_master_readdatavalid                          : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_data_master_readdatavalid -> nios2_gen2_0:d_readdatavalid
	signal nios2_gen2_0_data_master_write                                  : std_logic;                     -- nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	signal nios2_gen2_0_data_master_writedata                              : std_logic_vector(31 downto 0); -- nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	signal nios2_gen2_0_instruction_master_readdata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	signal nios2_gen2_0_instruction_master_waitrequest                     : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	signal nios2_gen2_0_instruction_master_address                         : std_logic_vector(20 downto 0); -- nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	signal nios2_gen2_0_instruction_master_read                            : std_logic;                     -- nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	signal nios2_gen2_0_instruction_master_readdatavalid                   : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_instruction_master_readdatavalid -> nios2_gen2_0:i_readdatavalid
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata         : std_logic_vector(31 downto 0); -- nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest      : std_logic;                     -- nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess      : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address          : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read             : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable       : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write            : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata        : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	signal mm_interconnect_0_sram_de2_0_s0_readdata                        : std_logic_vector(15 downto 0); -- SRAM_DE2_0:avs_s0_readdata -> mm_interconnect_0:SRAM_DE2_0_s0_readdata
	signal mm_interconnect_0_sram_de2_0_s0_address                         : std_logic_vector(17 downto 0); -- mm_interconnect_0:SRAM_DE2_0_s0_address -> SRAM_DE2_0:avs_s0_address
	signal mm_interconnect_0_sram_de2_0_s0_read                            : std_logic;                     -- mm_interconnect_0:SRAM_DE2_0_s0_read -> SRAM_DE2_0:avs_s0_read
	signal mm_interconnect_0_sram_de2_0_s0_byteenable                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:SRAM_DE2_0_s0_byteenable -> SRAM_DE2_0:avs_s0_byteenable
	signal mm_interconnect_0_sram_de2_0_s0_write                           : std_logic;                     -- mm_interconnect_0:SRAM_DE2_0_s0_write -> SRAM_DE2_0:avs_s0_write
	signal mm_interconnect_0_sram_de2_0_s0_writedata                       : std_logic_vector(15 downto 0); -- mm_interconnect_0:SRAM_DE2_0_s0_writedata -> SRAM_DE2_0:avs_s0_writedata
	signal mm_interconnect_0_pos_raquette_s1_readdata                      : std_logic_vector(31 downto 0); -- pos_raquette:readdata -> mm_interconnect_0:pos_raquette_s1_readdata
	signal mm_interconnect_0_pos_raquette_s1_address                       : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pos_raquette_s1_address -> pos_raquette:address
	signal mm_interconnect_0_brique_morte_s1_readdata                      : std_logic_vector(31 downto 0); -- brique_morte:readdata -> mm_interconnect_0:brique_morte_s1_readdata
	signal mm_interconnect_0_brique_morte_s1_address                       : std_logic_vector(1 downto 0);  -- mm_interconnect_0:brique_morte_s1_address -> brique_morte:address
	signal mm_interconnect_0_adr_brique_s1_chipselect                      : std_logic;                     -- mm_interconnect_0:adr_brique_s1_chipselect -> adr_brique:chipselect
	signal mm_interconnect_0_adr_brique_s1_readdata                        : std_logic_vector(31 downto 0); -- adr_brique:readdata -> mm_interconnect_0:adr_brique_s1_readdata
	signal mm_interconnect_0_adr_brique_s1_address                         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:adr_brique_s1_address -> adr_brique:address
	signal mm_interconnect_0_adr_brique_s1_write                           : std_logic;                     -- mm_interconnect_0:adr_brique_s1_write -> mm_interconnect_0_adr_brique_s1_write:in
	signal mm_interconnect_0_adr_brique_s1_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:adr_brique_s1_writedata -> adr_brique:writedata
	signal mm_interconnect_0_en_nios_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:en_nios_s1_chipselect -> en_nios:chipselect
	signal mm_interconnect_0_en_nios_s1_readdata                           : std_logic_vector(31 downto 0); -- en_nios:readdata -> mm_interconnect_0:en_nios_s1_readdata
	signal mm_interconnect_0_en_nios_s1_address                            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:en_nios_s1_address -> en_nios:address
	signal mm_interconnect_0_en_nios_s1_write                              : std_logic;                     -- mm_interconnect_0:en_nios_s1_write -> mm_interconnect_0_en_nios_s1_write:in
	signal mm_interconnect_0_en_nios_s1_writedata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:en_nios_s1_writedata -> en_nios:writedata
	signal mm_interconnect_0_perdu_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:perdu_s1_chipselect -> perdu:chipselect
	signal mm_interconnect_0_perdu_s1_readdata                             : std_logic_vector(31 downto 0); -- perdu:readdata -> mm_interconnect_0:perdu_s1_readdata
	signal mm_interconnect_0_perdu_s1_address                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:perdu_s1_address -> perdu:address
	signal mm_interconnect_0_perdu_s1_write                                : std_logic;                     -- mm_interconnect_0:perdu_s1_write -> mm_interconnect_0_perdu_s1_write:in
	signal mm_interconnect_0_perdu_s1_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:perdu_s1_writedata -> perdu:writedata
	signal mm_interconnect_0_en_s1_readdata                                : std_logic_vector(31 downto 0); -- en:readdata -> mm_interconnect_0:en_s1_readdata
	signal mm_interconnect_0_en_s1_address                                 : std_logic_vector(1 downto 0);  -- mm_interconnect_0:en_s1_address -> en:address
	signal mm_interconnect_0_fincalcul_s1_chipselect                       : std_logic;                     -- mm_interconnect_0:fincalcul_s1_chipselect -> fincalcul:chipselect
	signal mm_interconnect_0_fincalcul_s1_readdata                         : std_logic_vector(31 downto 0); -- fincalcul:readdata -> mm_interconnect_0:fincalcul_s1_readdata
	signal mm_interconnect_0_fincalcul_s1_address                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:fincalcul_s1_address -> fincalcul:address
	signal mm_interconnect_0_fincalcul_s1_write                            : std_logic;                     -- mm_interconnect_0:fincalcul_s1_write -> mm_interconnect_0_fincalcul_s1_write:in
	signal mm_interconnect_0_fincalcul_s1_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:fincalcul_s1_writedata -> fincalcul:writedata
	signal mm_interconnect_0_x_position_s1_chipselect                      : std_logic;                     -- mm_interconnect_0:x_position_s1_chipselect -> x_position:chipselect
	signal mm_interconnect_0_x_position_s1_readdata                        : std_logic_vector(31 downto 0); -- x_position:readdata -> mm_interconnect_0:x_position_s1_readdata
	signal mm_interconnect_0_x_position_s1_address                         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:x_position_s1_address -> x_position:address
	signal mm_interconnect_0_x_position_s1_write                           : std_logic;                     -- mm_interconnect_0:x_position_s1_write -> mm_interconnect_0_x_position_s1_write:in
	signal mm_interconnect_0_x_position_s1_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:x_position_s1_writedata -> x_position:writedata
	signal mm_interconnect_0_y_position_s1_chipselect                      : std_logic;                     -- mm_interconnect_0:y_position_s1_chipselect -> y_position:chipselect
	signal mm_interconnect_0_y_position_s1_readdata                        : std_logic_vector(31 downto 0); -- y_position:readdata -> mm_interconnect_0:y_position_s1_readdata
	signal mm_interconnect_0_y_position_s1_address                         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:y_position_s1_address -> y_position:address
	signal mm_interconnect_0_y_position_s1_write                           : std_logic;                     -- mm_interconnect_0:y_position_s1_write -> mm_interconnect_0_y_position_s1_write:in
	signal mm_interconnect_0_y_position_s1_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:y_position_s1_writedata -> y_position:writedata
	signal irq_mapper_receiver0_irq                                        : std_logic;                     -- jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	signal nios2_gen2_0_irq_irq                                            : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2_gen2_0:irq
	signal rst_controller_reset_out_reset                                  : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                              : std_logic;                     -- rst_controller:reset_req -> [nios2_gen2_0:reset_req, rst_translator:reset_req_in]
	signal nios2_gen2_0_debug_reset_request_reset                          : std_logic;                     -- nios2_gen2_0:debug_reset_request -> rst_controller:reset_in1
	signal reset_reset_n_ports_inv                                         : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:inv -> jtag_uart_0:av_read_n
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:inv -> jtag_uart_0:av_write_n
	signal mm_interconnect_0_adr_brique_s1_write_ports_inv                 : std_logic;                     -- mm_interconnect_0_adr_brique_s1_write:inv -> adr_brique:write_n
	signal mm_interconnect_0_en_nios_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_en_nios_s1_write:inv -> en_nios:write_n
	signal mm_interconnect_0_perdu_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_perdu_s1_write:inv -> perdu:write_n
	signal mm_interconnect_0_fincalcul_s1_write_ports_inv                  : std_logic;                     -- mm_interconnect_0_fincalcul_s1_write:inv -> fincalcul:write_n
	signal mm_interconnect_0_x_position_s1_write_ports_inv                 : std_logic;                     -- mm_interconnect_0_x_position_s1_write:inv -> x_position:write_n
	signal mm_interconnect_0_y_position_s1_write_ports_inv                 : std_logic;                     -- mm_interconnect_0_y_position_s1_write:inv -> y_position:write_n
	signal rst_controller_reset_out_reset_ports_inv                        : std_logic;                     -- rst_controller_reset_out_reset:inv -> [SRAM_DE2_0:reset_n, adr_brique:reset_n, brique_morte:reset_n, en:reset_n, en_nios:reset_n, fincalcul:reset_n, jtag_uart_0:rst_n, nios2_gen2_0:reset_n, perdu:reset_n, pos_raquette:reset_n, x_position:reset_n, y_position:reset_n]

begin

	sram_de2_0 : component SRAM_DE2
		port map (
			clk               => clk_clk,                                    --         clock.clk
			reset_n           => rst_controller_reset_out_reset_ports_inv,   --         reset.reset_n
			avs_s0_readdata   => mm_interconnect_0_sram_de2_0_s0_readdata,   --            s0.readdata
			avs_s0_writedata  => mm_interconnect_0_sram_de2_0_s0_writedata,  --              .writedata
			avs_s0_address    => mm_interconnect_0_sram_de2_0_s0_address,    --              .address
			avs_s0_write      => mm_interconnect_0_sram_de2_0_s0_write,      --              .write
			avs_s0_read       => mm_interconnect_0_sram_de2_0_s0_read,       --              .read
			avs_s0_byteenable => mm_interconnect_0_sram_de2_0_s0_byteenable, --              .byteenable
			coe_SRAM_ADDR     => sram_de2_ADDR,                              -- conduit_end_0.export
			coe_SRAM_DQ       => sram_de2_DQ,                                --              .export
			coe_SRAM_WE_N     => sram_de2_WE_N,                              --              .export
			coe_SRAM_OE_N     => sram_de2_OE_N,                              --              .export
			coe_SRAM_UB_N     => sram_de2_UB_N,                              --              .export
			coe_SRAM_LB_N     => sram_de2_LB_N,                              --              .export
			coe_SRAM_CE_N     => sram_de2_CE_N                               --              .export
		);

	adr_brique : component Niosballe_adr_brique
		port map (
			clk        => clk_clk,                                         --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,        --               reset.reset_n
			address    => mm_interconnect_0_adr_brique_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_adr_brique_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_adr_brique_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_adr_brique_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_adr_brique_s1_readdata,        --                    .readdata
			out_port   => adr_brique_export                                -- external_connection.export
		);

	brique_morte : component Niosballe_brique_morte
		port map (
			clk      => clk_clk,                                    --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address  => mm_interconnect_0_brique_morte_s1_address,  --                  s1.address
			readdata => mm_interconnect_0_brique_morte_s1_readdata, --                    .readdata
			in_port  => brique_morte_export                         -- external_connection.export
		);

	en : component Niosballe_brique_morte
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_en_s1_address,          --                  s1.address
			readdata => mm_interconnect_0_en_s1_readdata,         --                    .readdata
			in_port  => en_export                                 -- external_connection.export
		);

	en_nios : component Niosballe_en_nios
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_0_en_nios_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_en_nios_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_en_nios_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_en_nios_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_en_nios_s1_readdata,        --                    .readdata
			out_port   => en_nios_export                                -- external_connection.export
		);

	fincalcul : component Niosballe_en_nios
		port map (
			clk        => clk_clk,                                        --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,       --               reset.reset_n
			address    => mm_interconnect_0_fincalcul_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_fincalcul_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_fincalcul_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_fincalcul_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_fincalcul_s1_readdata,        --                    .readdata
			out_port   => fincalcul_export                                -- external_connection.export
		);

	jtag_uart_0 : component Niosballe_jtag_uart_0
		port map (
			clk            => clk_clk,                                                         --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                        --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                         --               irq.irq
		);

	nios2_gen2_0 : component Niosballe_nios2_gen2_0
		port map (
			clk                                 => clk_clk,                                                    --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,                   --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                         --                          .reset_req
			d_address                           => nios2_gen2_0_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_gen2_0_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_gen2_0_data_master_read,                              --                          .read
			d_readdata                          => nios2_gen2_0_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_gen2_0_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_gen2_0_data_master_write,                             --                          .write
			d_writedata                         => nios2_gen2_0_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => nios2_gen2_0_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => nios2_gen2_0_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_gen2_0_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_gen2_0_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_gen2_0_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_gen2_0_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => nios2_gen2_0_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => nios2_gen2_0_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios2_gen2_0_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                        -- custom_instruction_master.readra
		);

	perdu : component Niosballe_en_nios
		port map (
			clk        => clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_perdu_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_perdu_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_perdu_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_perdu_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_perdu_s1_readdata,        --                    .readdata
			out_port   => perdu_export                                -- external_connection.export
		);

	pos_raquette : component Niosballe_pos_raquette
		port map (
			clk      => clk_clk,                                    --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address  => mm_interconnect_0_pos_raquette_s1_address,  --                  s1.address
			readdata => mm_interconnect_0_pos_raquette_s1_readdata, --                    .readdata
			in_port  => pos_raquette_export                         -- external_connection.export
		);

	x_position : component Niosballe_x_position
		port map (
			clk        => clk_clk,                                         --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,        --               reset.reset_n
			address    => mm_interconnect_0_x_position_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_x_position_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_x_position_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_x_position_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_x_position_s1_readdata,        --                    .readdata
			out_port   => x_position_export                                -- external_connection.export
		);

	y_position : component Niosballe_x_position
		port map (
			clk        => clk_clk,                                         --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,        --               reset.reset_n
			address    => mm_interconnect_0_y_position_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_y_position_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_y_position_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_y_position_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_y_position_s1_readdata,        --                    .readdata
			out_port   => y_position_export                                -- external_connection.export
		);

	mm_interconnect_0 : component Niosballe_mm_interconnect_0
		port map (
			clk_0_clk_clk                                  => clk_clk,                                                     --                                clk_0_clk.clk
			nios2_gen2_0_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                              -- nios2_gen2_0_reset_reset_bridge_in_reset.reset
			nios2_gen2_0_data_master_address               => nios2_gen2_0_data_master_address,                            --                 nios2_gen2_0_data_master.address
			nios2_gen2_0_data_master_waitrequest           => nios2_gen2_0_data_master_waitrequest,                        --                                         .waitrequest
			nios2_gen2_0_data_master_byteenable            => nios2_gen2_0_data_master_byteenable,                         --                                         .byteenable
			nios2_gen2_0_data_master_read                  => nios2_gen2_0_data_master_read,                               --                                         .read
			nios2_gen2_0_data_master_readdata              => nios2_gen2_0_data_master_readdata,                           --                                         .readdata
			nios2_gen2_0_data_master_readdatavalid         => nios2_gen2_0_data_master_readdatavalid,                      --                                         .readdatavalid
			nios2_gen2_0_data_master_write                 => nios2_gen2_0_data_master_write,                              --                                         .write
			nios2_gen2_0_data_master_writedata             => nios2_gen2_0_data_master_writedata,                          --                                         .writedata
			nios2_gen2_0_data_master_debugaccess           => nios2_gen2_0_data_master_debugaccess,                        --                                         .debugaccess
			nios2_gen2_0_instruction_master_address        => nios2_gen2_0_instruction_master_address,                     --          nios2_gen2_0_instruction_master.address
			nios2_gen2_0_instruction_master_waitrequest    => nios2_gen2_0_instruction_master_waitrequest,                 --                                         .waitrequest
			nios2_gen2_0_instruction_master_read           => nios2_gen2_0_instruction_master_read,                        --                                         .read
			nios2_gen2_0_instruction_master_readdata       => nios2_gen2_0_instruction_master_readdata,                    --                                         .readdata
			nios2_gen2_0_instruction_master_readdatavalid  => nios2_gen2_0_instruction_master_readdatavalid,               --                                         .readdatavalid
			adr_brique_s1_address                          => mm_interconnect_0_adr_brique_s1_address,                     --                            adr_brique_s1.address
			adr_brique_s1_write                            => mm_interconnect_0_adr_brique_s1_write,                       --                                         .write
			adr_brique_s1_readdata                         => mm_interconnect_0_adr_brique_s1_readdata,                    --                                         .readdata
			adr_brique_s1_writedata                        => mm_interconnect_0_adr_brique_s1_writedata,                   --                                         .writedata
			adr_brique_s1_chipselect                       => mm_interconnect_0_adr_brique_s1_chipselect,                  --                                         .chipselect
			brique_morte_s1_address                        => mm_interconnect_0_brique_morte_s1_address,                   --                          brique_morte_s1.address
			brique_morte_s1_readdata                       => mm_interconnect_0_brique_morte_s1_readdata,                  --                                         .readdata
			en_s1_address                                  => mm_interconnect_0_en_s1_address,                             --                                    en_s1.address
			en_s1_readdata                                 => mm_interconnect_0_en_s1_readdata,                            --                                         .readdata
			en_nios_s1_address                             => mm_interconnect_0_en_nios_s1_address,                        --                               en_nios_s1.address
			en_nios_s1_write                               => mm_interconnect_0_en_nios_s1_write,                          --                                         .write
			en_nios_s1_readdata                            => mm_interconnect_0_en_nios_s1_readdata,                       --                                         .readdata
			en_nios_s1_writedata                           => mm_interconnect_0_en_nios_s1_writedata,                      --                                         .writedata
			en_nios_s1_chipselect                          => mm_interconnect_0_en_nios_s1_chipselect,                     --                                         .chipselect
			fincalcul_s1_address                           => mm_interconnect_0_fincalcul_s1_address,                      --                             fincalcul_s1.address
			fincalcul_s1_write                             => mm_interconnect_0_fincalcul_s1_write,                        --                                         .write
			fincalcul_s1_readdata                          => mm_interconnect_0_fincalcul_s1_readdata,                     --                                         .readdata
			fincalcul_s1_writedata                         => mm_interconnect_0_fincalcul_s1_writedata,                    --                                         .writedata
			fincalcul_s1_chipselect                        => mm_interconnect_0_fincalcul_s1_chipselect,                   --                                         .chipselect
			jtag_uart_0_avalon_jtag_slave_address          => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address,     --            jtag_uart_0_avalon_jtag_slave.address
			jtag_uart_0_avalon_jtag_slave_write            => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write,       --                                         .write
			jtag_uart_0_avalon_jtag_slave_read             => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read,        --                                         .read
			jtag_uart_0_avalon_jtag_slave_readdata         => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,    --                                         .readdata
			jtag_uart_0_avalon_jtag_slave_writedata        => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,   --                                         .writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest, --                                         .waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect       => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,  --                                         .chipselect
			nios2_gen2_0_debug_mem_slave_address           => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,      --             nios2_gen2_0_debug_mem_slave.address
			nios2_gen2_0_debug_mem_slave_write             => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,        --                                         .write
			nios2_gen2_0_debug_mem_slave_read              => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,         --                                         .read
			nios2_gen2_0_debug_mem_slave_readdata          => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,     --                                         .readdata
			nios2_gen2_0_debug_mem_slave_writedata         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,    --                                         .writedata
			nios2_gen2_0_debug_mem_slave_byteenable        => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,   --                                         .byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest       => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest,  --                                         .waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess       => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess,  --                                         .debugaccess
			perdu_s1_address                               => mm_interconnect_0_perdu_s1_address,                          --                                 perdu_s1.address
			perdu_s1_write                                 => mm_interconnect_0_perdu_s1_write,                            --                                         .write
			perdu_s1_readdata                              => mm_interconnect_0_perdu_s1_readdata,                         --                                         .readdata
			perdu_s1_writedata                             => mm_interconnect_0_perdu_s1_writedata,                        --                                         .writedata
			perdu_s1_chipselect                            => mm_interconnect_0_perdu_s1_chipselect,                       --                                         .chipselect
			pos_raquette_s1_address                        => mm_interconnect_0_pos_raquette_s1_address,                   --                          pos_raquette_s1.address
			pos_raquette_s1_readdata                       => mm_interconnect_0_pos_raquette_s1_readdata,                  --                                         .readdata
			SRAM_DE2_0_s0_address                          => mm_interconnect_0_sram_de2_0_s0_address,                     --                            SRAM_DE2_0_s0.address
			SRAM_DE2_0_s0_write                            => mm_interconnect_0_sram_de2_0_s0_write,                       --                                         .write
			SRAM_DE2_0_s0_read                             => mm_interconnect_0_sram_de2_0_s0_read,                        --                                         .read
			SRAM_DE2_0_s0_readdata                         => mm_interconnect_0_sram_de2_0_s0_readdata,                    --                                         .readdata
			SRAM_DE2_0_s0_writedata                        => mm_interconnect_0_sram_de2_0_s0_writedata,                   --                                         .writedata
			SRAM_DE2_0_s0_byteenable                       => mm_interconnect_0_sram_de2_0_s0_byteenable,                  --                                         .byteenable
			x_position_s1_address                          => mm_interconnect_0_x_position_s1_address,                     --                            x_position_s1.address
			x_position_s1_write                            => mm_interconnect_0_x_position_s1_write,                       --                                         .write
			x_position_s1_readdata                         => mm_interconnect_0_x_position_s1_readdata,                    --                                         .readdata
			x_position_s1_writedata                        => mm_interconnect_0_x_position_s1_writedata,                   --                                         .writedata
			x_position_s1_chipselect                       => mm_interconnect_0_x_position_s1_chipselect,                  --                                         .chipselect
			y_position_s1_address                          => mm_interconnect_0_y_position_s1_address,                     --                            y_position_s1.address
			y_position_s1_write                            => mm_interconnect_0_y_position_s1_write,                       --                                         .write
			y_position_s1_readdata                         => mm_interconnect_0_y_position_s1_readdata,                    --                                         .readdata
			y_position_s1_writedata                        => mm_interconnect_0_y_position_s1_writedata,                   --                                         .writedata
			y_position_s1_chipselect                       => mm_interconnect_0_y_position_s1_chipselect                   --                                         .chipselect
		);

	irq_mapper : component Niosballe_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			sender_irq    => nios2_gen2_0_irq_irq            --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                -- reset_in0.reset
			reset_in1      => nios2_gen2_0_debug_reset_request_reset, -- reset_in1.reset
			clk            => clk_clk,                                --       clk.clk
			reset_out      => rst_controller_reset_out_reset,         -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req,     --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;

	mm_interconnect_0_adr_brique_s1_write_ports_inv <= not mm_interconnect_0_adr_brique_s1_write;

	mm_interconnect_0_en_nios_s1_write_ports_inv <= not mm_interconnect_0_en_nios_s1_write;

	mm_interconnect_0_perdu_s1_write_ports_inv <= not mm_interconnect_0_perdu_s1_write;

	mm_interconnect_0_fincalcul_s1_write_ports_inv <= not mm_interconnect_0_fincalcul_s1_write;

	mm_interconnect_0_x_position_s1_write_ports_inv <= not mm_interconnect_0_x_position_s1_write;

	mm_interconnect_0_y_position_s1_write_ports_inv <= not mm_interconnect_0_y_position_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of Niosballe
